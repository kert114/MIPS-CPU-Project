module mips_cpu_bus_tb();
	