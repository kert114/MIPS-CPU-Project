module testfile(
	
);

	

endmodule :