module angus();
endmodule